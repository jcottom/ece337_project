module activation(
                  input wire [15:0]  in,
                  output wire [15:0] out
                  );
   reg [15:0]                       lut [0:65535] = '{
16'h00A4, 16'h00A4, 16'h00A4, 16'h00A5, 16'h00A5, 16'h00A5, 16'h00A5, 16'h00A6,
16'h00A6, 16'h00A6, 16'h00A6, 16'h00A7, 16'h00A7, 16'h00A7, 16'h00A7, 16'h00A8,
16'h00A8, 16'h00A8, 16'h00A8, 16'h00A9, 16'h00A9, 16'h00A9, 16'h00A9, 16'h00AA,
16'h00AA, 16'h00AA, 16'h00AA, 16'h00AB, 16'h00AB, 16'h00AB, 16'h00AB, 16'h00AC,
16'h00AC, 16'h00AC, 16'h00AC, 16'h00AD, 16'h00AD, 16'h00AD, 16'h00AD, 16'h00AE,
16'h00AE, 16'h00AE, 16'h00AE, 16'h00AF, 16'h00AF, 16'h00AF, 16'h00AF, 16'h00B0,
16'h00B0, 16'h00B0, 16'h00B0, 16'h00B1, 16'h00B1, 16'h00B1, 16'h00B1, 16'h00B2,
16'h00B2, 16'h00B2, 16'h00B2, 16'h00B3, 16'h00B3, 16'h00B3, 16'h00B3, 16'h00B4,
16'h00B4, 16'h00B4, 16'h00B4, 16'h00B5, 16'h00B5, 16'h00B5, 16'h00B5, 16'h00B6,
16'h00B6, 16'h00B6, 16'h00B6, 16'h00B7, 16'h00B7, 16'h00B7, 16'h00B7, 16'h00B7,
16'h00B8, 16'h00B8, 16'h00B8, 16'h00B8, 16'h00B9, 16'h00B9, 16'h00B9, 16'h00B9,
16'h00BA, 16'h00BA, 16'h00BA, 16'h00BA, 16'h00BB, 16'h00BB, 16'h00BB, 16'h00BB,
16'h00BC, 16'h00BC, 16'h00BC, 16'h00BC, 16'h00BD, 16'h00BD, 16'h00BD, 16'h00BD,
16'h00BE, 16'h00BE, 16'h00BE, 16'h00BE, 16'h00BF, 16'h00BF, 16'h00BF, 16'h00BF,
16'h00C0, 16'h00C0, 16'h00C0, 16'h00C0, 16'h00C1, 16'h00C1, 16'h00C1, 16'h00C1,
16'h00C2, 16'h00C2, 16'h00C2, 16'h00C2, 16'h00C2, 16'h00C3, 16'h00C3, 16'h00C3,
16'h00C3, 16'h00C4, 16'h00C4, 16'h00C4, 16'h00C4, 16'h00C5, 16'h00C5, 16'h00C5,
16'h00C5, 16'h00C6, 16'h00C6, 16'h00C6, 16'h00C6, 16'h00C7, 16'h00C7, 16'h00C7,
16'h00C7, 16'h00C8, 16'h00C8, 16'h00C8, 16'h00C8, 16'h00C8, 16'h00C9, 16'h00C9,
16'h00C9, 16'h00C9, 16'h00CA, 16'h00CA, 16'h00CA, 16'h00CA, 16'h00CB, 16'h00CB,
16'h00CB, 16'h00CB, 16'h00CC, 16'h00CC, 16'h00CC, 16'h00CC, 16'h00CC, 16'h00CD,
16'h00CD, 16'h00CD, 16'h00CD, 16'h00CE, 16'h00CE, 16'h00CE, 16'h00CE, 16'h00CF,
16'h00CF, 16'h00CF, 16'h00CF, 16'h00D0, 16'h00D0, 16'h00D0, 16'h00D0, 16'h00D0,
16'h00D1, 16'h00D1, 16'h00D1, 16'h00D1, 16'h00D2, 16'h00D2, 16'h00D2, 16'h00D2,
16'h00D3, 16'h00D3, 16'h00D3, 16'h00D3, 16'h00D3, 16'h00D4, 16'h00D4, 16'h00D4,
16'h00D4, 16'h00D5, 16'h00D5, 16'h00D5, 16'h00D5, 16'h00D5, 16'h00D6, 16'h00D6,
16'h00D6, 16'h00D6, 16'h00D7, 16'h00D7, 16'h00D7, 16'h00D7, 16'h00D8, 16'h00D8,
16'h00D8, 16'h00D8, 16'h00D8, 16'h00D9, 16'h00D9, 16'h00D9, 16'h00D9, 16'h00DA,
16'h00DA, 16'h00DA, 16'h00DA, 16'h00DA, 16'h00DB, 16'h00DB, 16'h00DB, 16'h00DB,
16'h00DC, 16'h00DC, 16'h00DC, 16'h00DC, 16'h00DC, 16'h00DD, 16'h00DD, 16'h00DD,
16'h00DD, 16'h00DE, 16'h00DE, 16'h00DE, 16'h00DE, 16'h00DE, 16'h00DF, 16'h00DF,
16'h00DF, 16'h00DF, 16'h00DF, 16'h00E0, 16'h00E0, 16'h00E0, 16'h00E0, 16'h00E1,
16'h00E1, 16'h00E1, 16'h00E1, 16'h00E1, 16'h00E2, 16'h00E2, 16'h00E2, 16'h00E2,
16'h00E2, 16'h00E3, 16'h00E3, 16'h00E3, 16'h00E3, 16'h00E4, 16'h00E4, 16'h00E4,
16'h00E4, 16'h00E4, 16'h00E5, 16'h00E5, 16'h00E5, 16'h00E5, 16'h00E5, 16'h00E6,
16'h00E6, 16'h00E6, 16'h00E6, 16'h00E6, 16'h00E7, 16'h00E7, 16'h00E7, 16'h00E7,
16'h00E8, 16'h00E8, 16'h00E8, 16'h00E8, 16'h00E8, 16'h00E9, 16'h00E9, 16'h00E9,
16'h00E9, 16'h00E9, 16'h00EA, 16'h00EA, 16'h00EA, 16'h00EA, 16'h00EA, 16'h00EB,
16'h00EB, 16'h00EB, 16'h00EB, 16'h00EB, 16'h00EC, 16'h00EC, 16'h00EC, 16'h00EC,
16'h00EC, 16'h00ED, 16'h00ED, 16'h00ED, 16'h00ED, 16'h00ED, 16'h00EE, 16'h00EE,
16'h00EE, 16'h00EE, 16'h00EE, 16'h00EF, 16'h00EF, 16'h00EF, 16'h00EF, 16'h00EF,
16'h00F0, 16'h00F0, 16'h00F0, 16'h00F0, 16'h00F0, 16'h00F1, 16'h00F1, 16'h00F1,
16'h00F1, 16'h00F1, 16'h00F2, 16'h00F2, 16'h00F2, 16'h00F2, 16'h00F2, 16'h00F3,
16'h00F3, 16'h00F3, 16'h00F3, 16'h00F3, 16'h00F3, 16'h00F4, 16'h00F4, 16'h00F4,
16'h00F4, 16'h00F4, 16'h00F5, 16'h00F5, 16'h00F5, 16'h00F5, 16'h00F5, 16'h00F6,
16'h00F6, 16'h00F6, 16'h00F6, 16'h00F6, 16'h00F7, 16'h00F7, 16'h00F7, 16'h00F7,
16'h00F7, 16'h00F7, 16'h00F8, 16'h00F8, 16'h00F8, 16'h00F8, 16'h00F8, 16'h00F9,
16'h00F9, 16'h00F9, 16'h00F9, 16'h00F9, 16'h00F9, 16'h00FA, 16'h00FA, 16'h00FA,
16'h00FA, 16'h00FA, 16'h00FB, 16'h00FB, 16'h00FB, 16'h00FB, 16'h00FB, 16'h00FB,
16'h00FC, 16'h00FC, 16'h00FC, 16'h00FC, 16'h00FC, 16'h00FC, 16'h00FD, 16'h00FD,
16'h00FD, 16'h00FD, 16'h00FD, 16'h00FE, 16'h00FE, 16'h00FE, 16'h00FE, 16'h00FE,
16'h00FE, 16'h00FF, 16'h00FF, 16'h00FF, 16'h00FF, 16'h00FF, 16'h00FF, 16'h0100,
16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0100, 16'h0101, 16'h0101, 16'h0101,
16'h0101, 16'h0101, 16'h0101, 16'h0102, 16'h0102, 16'h0102, 16'h0102, 16'h0102,
16'h0103, 16'h0103, 16'h0103, 16'h0103, 16'h0103, 16'h0103, 16'h0103, 16'h0104,
16'h0104, 16'h0104, 16'h0104, 16'h0104, 16'h0104, 16'h0105, 16'h0105, 16'h0105,
16'h0105, 16'h0105, 16'h0105, 16'h0106, 16'h0106, 16'h0106, 16'h0106, 16'h0106,
16'h0106, 16'h0107, 16'h0107, 16'h0107, 16'h0107, 16'h0107, 16'h0107, 16'h0108,
16'h0108, 16'h0108, 16'h0108, 16'h0108, 16'h0108, 16'h0108, 16'h0109, 16'h0109,
16'h0109, 16'h0109, 16'h0109, 16'h0109, 16'h010A, 16'h010A, 16'h010A, 16'h010A,
16'h010A, 16'h010A, 16'h010A, 16'h010B, 16'h010B, 16'h010B, 16'h010B, 16'h010B,
16'h010B, 16'h010C, 16'h010C, 16'h010C, 16'h010C, 16'h010C, 16'h010C, 16'h010C,
16'h010D, 16'h010D, 16'h010D, 16'h010D, 16'h010D, 16'h010D, 16'h010D, 16'h010E,
16'h010E, 16'h010E, 16'h010E, 16'h010E, 16'h010E, 16'h010E, 16'h010F, 16'h010F,
16'h010F, 16'h010F, 16'h010F, 16'h010F, 16'h010F, 16'h0110, 16'h0110, 16'h0110,
16'h0110, 16'h0110, 16'h0110, 16'h0110, 16'h0111, 16'h0111, 16'h0111, 16'h0111,
16'h0111, 16'h0111, 16'h0111, 16'h0112, 16'h0112, 16'h0112, 16'h0112, 16'h0112,
16'h0112, 16'h0112, 16'h0113, 16'h0113, 16'h0113, 16'h0113, 16'h0113, 16'h0113,
16'h0113, 16'h0113, 16'h0114, 16'h0114, 16'h0114, 16'h0114, 16'h0114, 16'h0114,
16'h0114, 16'h0115, 16'h0115, 16'h0115, 16'h0115, 16'h0115, 16'h0115, 16'h0115,
16'h0115, 16'h0116, 16'h0116, 16'h0116, 16'h0116, 16'h0116, 16'h0116, 16'h0116,
16'h0116, 16'h0117, 16'h0117, 16'h0117, 16'h0117, 16'h0117, 16'h0117, 16'h0117,
16'h0117, 16'h0118, 16'h0118, 16'h0118, 16'h0118, 16'h0118, 16'h0118, 16'h0118,
16'h0118, 16'h0119, 16'h0119, 16'h0119, 16'h0119, 16'h0119, 16'h0119, 16'h0119,
16'h0119, 16'h011A, 16'h011A, 16'h011A, 16'h011A, 16'h011A, 16'h011A, 16'h011A,
16'h011A, 16'h011B, 16'h011B, 16'h011B, 16'h011B, 16'h011B, 16'h011B, 16'h011B,
16'h011B, 16'h011B, 16'h011C, 16'h011C, 16'h011C, 16'h011C, 16'h011C, 16'h011C,
16'h011C, 16'h011C, 16'h011D, 16'h011D, 16'h011D, 16'h011D, 16'h011D, 16'h011D,
16'h011D, 16'h011D, 16'h011D, 16'h011E, 16'h011E, 16'h011E, 16'h011E, 16'h011E,
16'h011E, 16'h011E, 16'h011E, 16'h011E, 16'h011F, 16'h011F, 16'h011F, 16'h011F,
16'h011F, 16'h011F, 16'h011F, 16'h011F, 16'h011F, 16'h0120, 16'h0120, 16'h0120,
16'h0120, 16'h0120, 16'h0120, 16'h0120, 16'h0120, 16'h0120, 16'h0120, 16'h0121,
16'h0121, 16'h0121, 16'h0121, 16'h0121, 16'h0121, 16'h0121, 16'h0121, 16'h0121,
16'h0122, 16'h0122, 16'h0122, 16'h0122, 16'h0122, 16'h0122, 16'h0122, 16'h0122,
16'h0122, 16'h0122, 16'h0123, 16'h0123, 16'h0123, 16'h0123, 16'h0123, 16'h0123,
16'h0123, 16'h0123, 16'h0123, 16'h0123, 16'h0124, 16'h0124, 16'h0124, 16'h0124,
16'h0124, 16'h0124, 16'h0124, 16'h0124, 16'h0124, 16'h0124, 16'h0124, 16'h0125,
16'h0125, 16'h0125, 16'h0125, 16'h0125, 16'h0125, 16'h0125, 16'h0125, 16'h0125,
16'h0125, 16'h0126, 16'h0126, 16'h0126, 16'h0126, 16'h0126, 16'h0126, 16'h0126,
16'h0126, 16'h0126, 16'h0126, 16'h0126, 16'h0127, 16'h0127, 16'h0127, 16'h0127,
16'h0127, 16'h0127, 16'h0127, 16'h0127, 16'h0127, 16'h0127, 16'h0127, 16'h0128,
16'h0128, 16'h0128, 16'h0128, 16'h0128, 16'h0128, 16'h0128, 16'h0128, 16'h0128,
16'h0128, 16'h0128, 16'h0128, 16'h0129, 16'h0129, 16'h0129, 16'h0129, 16'h0129,
16'h0129, 16'h0129, 16'h0129, 16'h0129, 16'h0129, 16'h0129, 16'h012A, 16'h012A,
16'h012A, 16'h012A, 16'h012A, 16'h012A, 16'h012A, 16'h012A, 16'h012A, 16'h012A,
16'h012A, 16'h012A, 16'h012A, 16'h012B, 16'h012B, 16'h012B, 16'h012B, 16'h012B,
16'h012B, 16'h012B, 16'h012B, 16'h012B, 16'h012B, 16'h012B, 16'h012B, 16'h012C,
16'h012C, 16'h012C, 16'h012C, 16'h012C, 16'h012C, 16'h012C, 16'h012C, 16'h012C,
16'h012C, 16'h012C, 16'h012C, 16'h012C, 16'h012D, 16'h012D, 16'h012D, 16'h012D,
16'h012D, 16'h012D, 16'h012D, 16'h012D, 16'h012D, 16'h012D, 16'h012D, 16'h012D,
16'h012D, 16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012E,
16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012E, 16'h012F,
16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h012F,
16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h012F, 16'h0130, 16'h0130,
16'h0130, 16'h0130, 16'h0130, 16'h0130, 16'h0130, 16'h0130, 16'h0130, 16'h0130,
16'h0130, 16'h0130, 16'h0130, 16'h0130, 16'h0130, 16'h0131, 16'h0131, 16'h0131,
16'h0131, 16'h0131, 16'h0131, 16'h0131, 16'h0131, 16'h0131, 16'h0131, 16'h0131,
16'h0131, 16'h0131, 16'h0131, 16'h0131, 16'h0132, 16'h0132, 16'h0132, 16'h0132,
16'h0132, 16'h0132, 16'h0132, 16'h0132, 16'h0132, 16'h0132, 16'h0132, 16'h0132,
16'h0132, 16'h0132, 16'h0132, 16'h0132, 16'h0133, 16'h0133, 16'h0133, 16'h0133,
16'h0133, 16'h0133, 16'h0133, 16'h0133, 16'h0133, 16'h0133, 16'h0133, 16'h0133,
16'h0133, 16'h0133, 16'h0133, 16'h0133, 16'h0133, 16'h0134, 16'h0134, 16'h0134,
16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134,
16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0134, 16'h0135,
16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135,
16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135, 16'h0135,
16'h0135, 16'h0135, 16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136,
16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136,
16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0136, 16'h0137, 16'h0137, 16'h0137,
16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137,
16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137, 16'h0137,
16'h0137, 16'h0137, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138,
16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138,
16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138, 16'h0138,
16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139,
16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139,
16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h0139, 16'h013A,
16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A,
16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A,
16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A, 16'h013A,
16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B,
16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B,
16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B, 16'h013B,
16'h013B, 16'h013B, 16'h013B, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C,
16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C,
16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C,
16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C, 16'h013C,
16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D,
16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D,
16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D,
16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D, 16'h013D,
16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E,
16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E,
16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E,
16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E, 16'h013E,
16'h013E, 16'h013E, 16'h013E, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F,
16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F,
16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F,
16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F,
16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F, 16'h013F,
16'h013F, 16'h013F, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140,
16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140,
16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140,
16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140,
16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140,
16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0140, 16'h0141, 16'h0141,
16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141,
16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141,
16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141,
16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141,
16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141,
16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141, 16'h0141,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142, 16'h0142,
16'h0142, 16'h0142, 16'h0142, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143, 16'h0143,
16'h0143, 16'h0143, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144,
16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0144, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145, 16'h0145,
16'h0145, 16'h0145, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146,
16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0146, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147,
16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0147, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148, 16'h0148,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000B, 16'h000B, 16'h000B, 16'h000B,
16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B,
16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B,
16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B,
16'h000B, 16'h000B, 16'h000B, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C,
16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C,
16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C,
16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000D,
16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D,
16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D,
16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D,
16'h000D, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E,
16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E,
16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E,
16'h000E, 16'h000E, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F,
16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F,
16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F,
16'h000F, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010,
16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010,
16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0011, 16'h0011,
16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011,
16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011,
16'h0011, 16'h0011, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012,
16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012,
16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0013, 16'h0013,
16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013,
16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013,
16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014,
16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014,
16'h0014, 16'h0014, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015,
16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015,
16'h0015, 16'h0015, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016,
16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016,
16'h0016, 16'h0016, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017,
16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017,
16'h0017, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018,
16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018,
16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019,
16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h001A, 16'h001A,
16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A,
16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001B, 16'h001B, 16'h001B, 16'h001B,
16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B,
16'h001B, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C,
16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001D, 16'h001D,
16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001D,
16'h001D, 16'h001D, 16'h001D, 16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001E,
16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001F,
16'h001F, 16'h001F, 16'h001F, 16'h001F, 16'h001F, 16'h001F, 16'h001F, 16'h001F,
16'h001F, 16'h001F, 16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0020,
16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0021, 16'h0021,
16'h0021, 16'h0021, 16'h0021, 16'h0021, 16'h0021, 16'h0021, 16'h0021, 16'h0021,
16'h0021, 16'h0022, 16'h0022, 16'h0022, 16'h0022, 16'h0022, 16'h0022, 16'h0022,
16'h0022, 16'h0022, 16'h0022, 16'h0023, 16'h0023, 16'h0023, 16'h0023, 16'h0023,
16'h0023, 16'h0023, 16'h0023, 16'h0023, 16'h0023, 16'h0023, 16'h0024, 16'h0024,
16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0024,
16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025,
16'h0025, 16'h0025, 16'h0026, 16'h0026, 16'h0026, 16'h0026, 16'h0026, 16'h0026,
16'h0026, 16'h0026, 16'h0026, 16'h0026, 16'h0027, 16'h0027, 16'h0027, 16'h0027,
16'h0027, 16'h0027, 16'h0027, 16'h0027, 16'h0027, 16'h0028, 16'h0028, 16'h0028,
16'h0028, 16'h0028, 16'h0028, 16'h0028, 16'h0028, 16'h0028, 16'h0028, 16'h0029,
16'h0029, 16'h0029, 16'h0029, 16'h0029, 16'h0029, 16'h0029, 16'h0029, 16'h0029,
16'h002A, 16'h002A, 16'h002A, 16'h002A, 16'h002A, 16'h002A, 16'h002A, 16'h002A,
16'h002A, 16'h002B, 16'h002B, 16'h002B, 16'h002B, 16'h002B, 16'h002B, 16'h002B,
16'h002B, 16'h002B, 16'h002C, 16'h002C, 16'h002C, 16'h002C, 16'h002C, 16'h002C,
16'h002C, 16'h002C, 16'h002D, 16'h002D, 16'h002D, 16'h002D, 16'h002D, 16'h002D,
16'h002D, 16'h002D, 16'h002D, 16'h002E, 16'h002E, 16'h002E, 16'h002E, 16'h002E,
16'h002E, 16'h002E, 16'h002E, 16'h002F, 16'h002F, 16'h002F, 16'h002F, 16'h002F,
16'h002F, 16'h002F, 16'h002F, 16'h0030, 16'h0030, 16'h0030, 16'h0030, 16'h0030,
16'h0030, 16'h0030, 16'h0030, 16'h0031, 16'h0031, 16'h0031, 16'h0031, 16'h0031,
16'h0031, 16'h0031, 16'h0031, 16'h0032, 16'h0032, 16'h0032, 16'h0032, 16'h0032,
16'h0032, 16'h0032, 16'h0032, 16'h0033, 16'h0033, 16'h0033, 16'h0033, 16'h0033,
16'h0033, 16'h0033, 16'h0034, 16'h0034, 16'h0034, 16'h0034, 16'h0034, 16'h0034,
16'h0034, 16'h0034, 16'h0035, 16'h0035, 16'h0035, 16'h0035, 16'h0035, 16'h0035,
16'h0035, 16'h0036, 16'h0036, 16'h0036, 16'h0036, 16'h0036, 16'h0036, 16'h0036,
16'h0037, 16'h0037, 16'h0037, 16'h0037, 16'h0037, 16'h0037, 16'h0037, 16'h0038,
16'h0038, 16'h0038, 16'h0038, 16'h0038, 16'h0038, 16'h0038, 16'h0038, 16'h0039,
16'h0039, 16'h0039, 16'h0039, 16'h0039, 16'h0039, 16'h0039, 16'h003A, 16'h003A,
16'h003A, 16'h003A, 16'h003A, 16'h003A, 16'h003B, 16'h003B, 16'h003B, 16'h003B,
16'h003B, 16'h003B, 16'h003B, 16'h003C, 16'h003C, 16'h003C, 16'h003C, 16'h003C,
16'h003C, 16'h003C, 16'h003D, 16'h003D, 16'h003D, 16'h003D, 16'h003D, 16'h003D,
16'h003E, 16'h003E, 16'h003E, 16'h003E, 16'h003E, 16'h003E, 16'h003E, 16'h003F,
16'h003F, 16'h003F, 16'h003F, 16'h003F, 16'h003F, 16'h0040, 16'h0040, 16'h0040,
16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0041, 16'h0041, 16'h0041, 16'h0041,
16'h0041, 16'h0041, 16'h0042, 16'h0042, 16'h0042, 16'h0042, 16'h0042, 16'h0042,
16'h0043, 16'h0043, 16'h0043, 16'h0043, 16'h0043, 16'h0043, 16'h0044, 16'h0044,
16'h0044, 16'h0044, 16'h0044, 16'h0044, 16'h0045, 16'h0045, 16'h0045, 16'h0045,
16'h0045, 16'h0045, 16'h0045, 16'h0046, 16'h0046, 16'h0046, 16'h0046, 16'h0046,
16'h0047, 16'h0047, 16'h0047, 16'h0047, 16'h0047, 16'h0047, 16'h0048, 16'h0048,
16'h0048, 16'h0048, 16'h0048, 16'h0048, 16'h0049, 16'h0049, 16'h0049, 16'h0049,
16'h0049, 16'h0049, 16'h004A, 16'h004A, 16'h004A, 16'h004A, 16'h004A, 16'h004A,
16'h004B, 16'h004B, 16'h004B, 16'h004B, 16'h004B, 16'h004C, 16'h004C, 16'h004C,
16'h004C, 16'h004C, 16'h004C, 16'h004D, 16'h004D, 16'h004D, 16'h004D, 16'h004D,
16'h004D, 16'h004E, 16'h004E, 16'h004E, 16'h004E, 16'h004E, 16'h004F, 16'h004F,
16'h004F, 16'h004F, 16'h004F, 16'h0050, 16'h0050, 16'h0050, 16'h0050, 16'h0050,
16'h0050, 16'h0051, 16'h0051, 16'h0051, 16'h0051, 16'h0051, 16'h0052, 16'h0052,
16'h0052, 16'h0052, 16'h0052, 16'h0052, 16'h0053, 16'h0053, 16'h0053, 16'h0053,
16'h0053, 16'h0054, 16'h0054, 16'h0054, 16'h0054, 16'h0054, 16'h0055, 16'h0055,
16'h0055, 16'h0055, 16'h0055, 16'h0056, 16'h0056, 16'h0056, 16'h0056, 16'h0056,
16'h0056, 16'h0057, 16'h0057, 16'h0057, 16'h0057, 16'h0057, 16'h0058, 16'h0058,
16'h0058, 16'h0058, 16'h0058, 16'h0059, 16'h0059, 16'h0059, 16'h0059, 16'h0059,
16'h005A, 16'h005A, 16'h005A, 16'h005A, 16'h005A, 16'h005B, 16'h005B, 16'h005B,
16'h005B, 16'h005B, 16'h005C, 16'h005C, 16'h005C, 16'h005C, 16'h005C, 16'h005D,
16'h005D, 16'h005D, 16'h005D, 16'h005D, 16'h005E, 16'h005E, 16'h005E, 16'h005E,
16'h005E, 16'h005F, 16'h005F, 16'h005F, 16'h005F, 16'h0060, 16'h0060, 16'h0060,
16'h0060, 16'h0060, 16'h0061, 16'h0061, 16'h0061, 16'h0061, 16'h0061, 16'h0062,
16'h0062, 16'h0062, 16'h0062, 16'h0062, 16'h0063, 16'h0063, 16'h0063, 16'h0063,
16'h0063, 16'h0064, 16'h0064, 16'h0064, 16'h0064, 16'h0065, 16'h0065, 16'h0065,
16'h0065, 16'h0065, 16'h0066, 16'h0066, 16'h0066, 16'h0066, 16'h0066, 16'h0067,
16'h0067, 16'h0067, 16'h0067, 16'h0068, 16'h0068, 16'h0068, 16'h0068, 16'h0068,
16'h0069, 16'h0069, 16'h0069, 16'h0069, 16'h006A, 16'h006A, 16'h006A, 16'h006A,
16'h006A, 16'h006B, 16'h006B, 16'h006B, 16'h006B, 16'h006B, 16'h006C, 16'h006C,
16'h006C, 16'h006C, 16'h006D, 16'h006D, 16'h006D, 16'h006D, 16'h006D, 16'h006E,
16'h006E, 16'h006E, 16'h006E, 16'h006F, 16'h006F, 16'h006F, 16'h006F, 16'h006F,
16'h0070, 16'h0070, 16'h0070, 16'h0070, 16'h0071, 16'h0071, 16'h0071, 16'h0071,
16'h0072, 16'h0072, 16'h0072, 16'h0072, 16'h0072, 16'h0073, 16'h0073, 16'h0073,
16'h0073, 16'h0074, 16'h0074, 16'h0074, 16'h0074, 16'h0074, 16'h0075, 16'h0075,
16'h0075, 16'h0075, 16'h0076, 16'h0076, 16'h0076, 16'h0076, 16'h0077, 16'h0077,
16'h0077, 16'h0077, 16'h0077, 16'h0078, 16'h0078, 16'h0078, 16'h0078, 16'h0079,
16'h0079, 16'h0079, 16'h0079, 16'h007A, 16'h007A, 16'h007A, 16'h007A, 16'h007A,
16'h007B, 16'h007B, 16'h007B, 16'h007B, 16'h007C, 16'h007C, 16'h007C, 16'h007C,
16'h007D, 16'h007D, 16'h007D, 16'h007D, 16'h007E, 16'h007E, 16'h007E, 16'h007E,
16'h007F, 16'h007F, 16'h007F, 16'h007F, 16'h007F, 16'h0080, 16'h0080, 16'h0080,
16'h0080, 16'h0081, 16'h0081, 16'h0081, 16'h0081, 16'h0082, 16'h0082, 16'h0082,
16'h0082, 16'h0083, 16'h0083, 16'h0083, 16'h0083, 16'h0084, 16'h0084, 16'h0084,
16'h0084, 16'h0084, 16'h0085, 16'h0085, 16'h0085, 16'h0085, 16'h0086, 16'h0086,
16'h0086, 16'h0086, 16'h0087, 16'h0087, 16'h0087, 16'h0087, 16'h0088, 16'h0088,
16'h0088, 16'h0088, 16'h0089, 16'h0089, 16'h0089, 16'h0089, 16'h008A, 16'h008A,
16'h008A, 16'h008A, 16'h008B, 16'h008B, 16'h008B, 16'h008B, 16'h008C, 16'h008C,
16'h008C, 16'h008C, 16'h008C, 16'h008D, 16'h008D, 16'h008D, 16'h008D, 16'h008E,
16'h008E, 16'h008E, 16'h008E, 16'h008F, 16'h008F, 16'h008F, 16'h008F, 16'h0090,
16'h0090, 16'h0090, 16'h0090, 16'h0091, 16'h0091, 16'h0091, 16'h0091, 16'h0092,
16'h0092, 16'h0092, 16'h0092, 16'h0093, 16'h0093, 16'h0093, 16'h0093, 16'h0094,
16'h0094, 16'h0094, 16'h0094, 16'h0095, 16'h0095, 16'h0095, 16'h0095, 16'h0096,
16'h0096, 16'h0096, 16'h0096, 16'h0097, 16'h0097, 16'h0097, 16'h0097, 16'h0098,
16'h0098, 16'h0098, 16'h0098, 16'h0099, 16'h0099, 16'h0099, 16'h0099, 16'h009A,
16'h009A, 16'h009A, 16'h009A, 16'h009B, 16'h009B, 16'h009B, 16'h009B, 16'h009C,
16'h009C, 16'h009C, 16'h009C, 16'h009D, 16'h009D, 16'h009D, 16'h009D, 16'h009E,
16'h009E, 16'h009E, 16'h009E, 16'h009F, 16'h009F, 16'h009F, 16'h009F, 16'h00A0,
16'h00A0, 16'h00A0, 16'h00A0, 16'h00A1, 16'h00A1, 16'h00A1, 16'h00A1, 16'h00A2,
16'h00A2, 16'h00A2, 16'h00A2, 16'h00A3, 16'h00A3, 16'h00A3, 16'h00A3, 16'h00A4
                                                      };
   assign out = lut[in];

endmodule // activation
