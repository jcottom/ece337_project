module read_file();


endmodule
