// $Id: $
// File name:   controller.sv
// Created:     11/8/2016
// Author:      Cheyenne Martinez
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: ANN Controller
