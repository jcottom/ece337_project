/*
 This module serves as the activation function for the neural network.  It is a
 combinational block which implements a look-up table for the sigmoid function:

                            f(x) = (1 + e^-x)^-1

 I assume that this table is synthesized as a 2^16 to 1 multiplexer, or a
 2^16*16 bit to 1*16 bit mux, which can be implemented as the following number
 of NAND gates:

      16*4(2^16/2 + 2^15/2 + ... + 2^2/2 + 2/2) = 16*4(2^16 - 1) = 4194240

 The current table entries assume a fixed-point encoding of

                      (0111 1111 1111 1111)_2 = 100_10
                      (0000 0000 0000 0000)_2 = 0_10

 This can be changed as needed by generating a new set of table entries with the
 script in ece337_project/python/lut.py. The variable s contains the scaling
 factor for the fixed point encoding, and the function genLUTArray() will print
 a new set of values for this table.  In order to test this design, one would
 need to generate a new ece337_project/python/lut.pat using the same scaling
 factor, which is used by the tb_activation module.
 */
module activation(
                  input wire [15:0]  in,
                  output wire [15:0] out
                  );
   reg [15:0]                       lut [0:65535] = '{
16'h0800, 16'h0804, 16'h0808, 16'h080C, 16'h0810, 16'h0814, 16'h0818, 16'h081C,
16'h0820, 16'h0824, 16'h0828, 16'h082C, 16'h0830, 16'h0834, 16'h0838, 16'h083C,
16'h0840, 16'h0844, 16'h0848, 16'h084C, 16'h0850, 16'h0854, 16'h0858, 16'h085C,
16'h0860, 16'h0864, 16'h0868, 16'h086C, 16'h0870, 16'h0874, 16'h0878, 16'h087C,
16'h0880, 16'h0884, 16'h0888, 16'h088C, 16'h0890, 16'h0894, 16'h0898, 16'h089C,
16'h08A0, 16'h08A4, 16'h08A8, 16'h08AC, 16'h08B0, 16'h08B4, 16'h08B8, 16'h08BB,
16'h08BF, 16'h08C3, 16'h08C7, 16'h08CB, 16'h08CF, 16'h08D3, 16'h08D7, 16'h08DB,
16'h08DF, 16'h08E3, 16'h08E7, 16'h08EB, 16'h08EF, 16'h08F3, 16'h08F7, 16'h08FB,
16'h08FF, 16'h0903, 16'h0907, 16'h090A, 16'h090E, 16'h0912, 16'h0916, 16'h091A,
16'h091E, 16'h0922, 16'h0926, 16'h092A, 16'h092E, 16'h0932, 16'h0936, 16'h093A,
16'h093D, 16'h0941, 16'h0945, 16'h0949, 16'h094D, 16'h0951, 16'h0955, 16'h0959,
16'h095D, 16'h0960, 16'h0964, 16'h0968, 16'h096C, 16'h0970, 16'h0974, 16'h0978,
16'h097C, 16'h097F, 16'h0983, 16'h0987, 16'h098B, 16'h098F, 16'h0993, 16'h0997,
16'h099A, 16'h099E, 16'h09A2, 16'h09A6, 16'h09AA, 16'h09AE, 16'h09B1, 16'h09B5,
16'h09B9, 16'h09BD, 16'h09C1, 16'h09C4, 16'h09C8, 16'h09CC, 16'h09D0, 16'h09D4,
16'h09D7, 16'h09DB, 16'h09DF, 16'h09E3, 16'h09E7, 16'h09EA, 16'h09EE, 16'h09F2,
16'h09F6, 16'h09F9, 16'h09FD, 16'h0A01, 16'h0A05, 16'h0A08, 16'h0A0C, 16'h0A10,
16'h0A14, 16'h0A17, 16'h0A1B, 16'h0A1F, 16'h0A22, 16'h0A26, 16'h0A2A, 16'h0A2E,
16'h0A31, 16'h0A35, 16'h0A39, 16'h0A3C, 16'h0A40, 16'h0A44, 16'h0A47, 16'h0A4B,
16'h0A4F, 16'h0A52, 16'h0A56, 16'h0A5A, 16'h0A5D, 16'h0A61, 16'h0A65, 16'h0A68,
16'h0A6C, 16'h0A70, 16'h0A73, 16'h0A77, 16'h0A7A, 16'h0A7E, 16'h0A82, 16'h0A85,
16'h0A89, 16'h0A8C, 16'h0A90, 16'h0A94, 16'h0A97, 16'h0A9B, 16'h0A9E, 16'h0AA2,
16'h0AA6, 16'h0AA9, 16'h0AAD, 16'h0AB0, 16'h0AB4, 16'h0AB7, 16'h0ABB, 16'h0ABE,
16'h0AC2, 16'h0AC5, 16'h0AC9, 16'h0ACC, 16'h0AD0, 16'h0AD3, 16'h0AD7, 16'h0ADA,
16'h0ADE, 16'h0AE1, 16'h0AE5, 16'h0AE8, 16'h0AEC, 16'h0AEF, 16'h0AF3, 16'h0AF6,
16'h0AFA, 16'h0AFD, 16'h0B01, 16'h0B04, 16'h0B07, 16'h0B0B, 16'h0B0E, 16'h0B12,
16'h0B15, 16'h0B18, 16'h0B1C, 16'h0B1F, 16'h0B23, 16'h0B26, 16'h0B29, 16'h0B2D,
16'h0B30, 16'h0B34, 16'h0B37, 16'h0B3A, 16'h0B3E, 16'h0B41, 16'h0B44, 16'h0B48,
16'h0B4B, 16'h0B4E, 16'h0B52, 16'h0B55, 16'h0B58, 16'h0B5B, 16'h0B5F, 16'h0B62,
16'h0B65, 16'h0B69, 16'h0B6C, 16'h0B6F, 16'h0B72, 16'h0B76, 16'h0B79, 16'h0B7C,
16'h0B7F, 16'h0B83, 16'h0B86, 16'h0B89, 16'h0B8C, 16'h0B8F, 16'h0B93, 16'h0B96,
16'h0B99, 16'h0B9C, 16'h0B9F, 16'h0BA3, 16'h0BA6, 16'h0BA9, 16'h0BAC, 16'h0BAF,
16'h0BB2, 16'h0BB6, 16'h0BB9, 16'h0BBC, 16'h0BBF, 16'h0BC2, 16'h0BC5, 16'h0BC8,
16'h0BCB, 16'h0BCE, 16'h0BD2, 16'h0BD5, 16'h0BD8, 16'h0BDB, 16'h0BDE, 16'h0BE1,
16'h0BE4, 16'h0BE7, 16'h0BEA, 16'h0BED, 16'h0BF0, 16'h0BF3, 16'h0BF6, 16'h0BF9,
16'h0BFC, 16'h0BFF, 16'h0C02, 16'h0C05, 16'h0C08, 16'h0C0B, 16'h0C0E, 16'h0C11,
16'h0C14, 16'h0C17, 16'h0C1A, 16'h0C1D, 16'h0C20, 16'h0C23, 16'h0C26, 16'h0C29,
16'h0C2C, 16'h0C2F, 16'h0C31, 16'h0C34, 16'h0C37, 16'h0C3A, 16'h0C3D, 16'h0C40,
16'h0C43, 16'h0C46, 16'h0C48, 16'h0C4B, 16'h0C4E, 16'h0C51, 16'h0C54, 16'h0C57,
16'h0C59, 16'h0C5C, 16'h0C5F, 16'h0C62, 16'h0C65, 16'h0C67, 16'h0C6A, 16'h0C6D,
16'h0C70, 16'h0C73, 16'h0C75, 16'h0C78, 16'h0C7B, 16'h0C7E, 16'h0C80, 16'h0C83,
16'h0C86, 16'h0C89, 16'h0C8B, 16'h0C8E, 16'h0C91, 16'h0C93, 16'h0C96, 16'h0C99,
16'h0C9B, 16'h0C9E, 16'h0CA1, 16'h0CA3, 16'h0CA6, 16'h0CA9, 16'h0CAB, 16'h0CAE,
16'h0CB1, 16'h0CB3, 16'h0CB6, 16'h0CB8, 16'h0CBB, 16'h0CBE, 16'h0CC0, 16'h0CC3,
16'h0CC5, 16'h0CC8, 16'h0CCB, 16'h0CCD, 16'h0CD0, 16'h0CD2, 16'h0CD5, 16'h0CD7,
16'h0CDA, 16'h0CDC, 16'h0CDF, 16'h0CE1, 16'h0CE4, 16'h0CE6, 16'h0CE9, 16'h0CEB,
16'h0CEE, 16'h0CF0, 16'h0CF3, 16'h0CF5, 16'h0CF8, 16'h0CFA, 16'h0CFD, 16'h0CFF,
16'h0D02, 16'h0D04, 16'h0D06, 16'h0D09, 16'h0D0B, 16'h0D0E, 16'h0D10, 16'h0D12,
16'h0D15, 16'h0D17, 16'h0D1A, 16'h0D1C, 16'h0D1E, 16'h0D21, 16'h0D23, 16'h0D25,
16'h0D28, 16'h0D2A, 16'h0D2C, 16'h0D2F, 16'h0D31, 16'h0D33, 16'h0D36, 16'h0D38,
16'h0D3A, 16'h0D3D, 16'h0D3F, 16'h0D41, 16'h0D43, 16'h0D46, 16'h0D48, 16'h0D4A,
16'h0D4C, 16'h0D4F, 16'h0D51, 16'h0D53, 16'h0D55, 16'h0D58, 16'h0D5A, 16'h0D5C,
16'h0D5E, 16'h0D60, 16'h0D63, 16'h0D65, 16'h0D67, 16'h0D69, 16'h0D6B, 16'h0D6D,
16'h0D70, 16'h0D72, 16'h0D74, 16'h0D76, 16'h0D78, 16'h0D7A, 16'h0D7C, 16'h0D7E,
16'h0D81, 16'h0D83, 16'h0D85, 16'h0D87, 16'h0D89, 16'h0D8B, 16'h0D8D, 16'h0D8F,
16'h0D91, 16'h0D93, 16'h0D95, 16'h0D97, 16'h0D99, 16'h0D9C, 16'h0D9E, 16'h0DA0,
16'h0DA2, 16'h0DA4, 16'h0DA6, 16'h0DA8, 16'h0DAA, 16'h0DAC, 16'h0DAE, 16'h0DB0,
16'h0DB2, 16'h0DB4, 16'h0DB6, 16'h0DB7, 16'h0DB9, 16'h0DBB, 16'h0DBD, 16'h0DBF,
16'h0DC1, 16'h0DC3, 16'h0DC5, 16'h0DC7, 16'h0DC9, 16'h0DCB, 16'h0DCD, 16'h0DCF,
16'h0DD0, 16'h0DD2, 16'h0DD4, 16'h0DD6, 16'h0DD8, 16'h0DDA, 16'h0DDC, 16'h0DDE,
16'h0DDF, 16'h0DE1, 16'h0DE3, 16'h0DE5, 16'h0DE7, 16'h0DE9, 16'h0DEA, 16'h0DEC,
16'h0DEE, 16'h0DF0, 16'h0DF2, 16'h0DF3, 16'h0DF5, 16'h0DF7, 16'h0DF9, 16'h0DFA,
16'h0DFC, 16'h0DFE, 16'h0E00, 16'h0E01, 16'h0E03, 16'h0E05, 16'h0E07, 16'h0E08,
16'h0E0A, 16'h0E0C, 16'h0E0E, 16'h0E0F, 16'h0E11, 16'h0E13, 16'h0E14, 16'h0E16,
16'h0E18, 16'h0E19, 16'h0E1B, 16'h0E1D, 16'h0E1E, 16'h0E20, 16'h0E22, 16'h0E23,
16'h0E25, 16'h0E27, 16'h0E28, 16'h0E2A, 16'h0E2C, 16'h0E2D, 16'h0E2F, 16'h0E30,
16'h0E32, 16'h0E34, 16'h0E35, 16'h0E37, 16'h0E38, 16'h0E3A, 16'h0E3C, 16'h0E3D,
16'h0E3F, 16'h0E40, 16'h0E42, 16'h0E43, 16'h0E45, 16'h0E46, 16'h0E48, 16'h0E49,
16'h0E4B, 16'h0E4D, 16'h0E4E, 16'h0E50, 16'h0E51, 16'h0E53, 16'h0E54, 16'h0E56,
16'h0E57, 16'h0E59, 16'h0E5A, 16'h0E5B, 16'h0E5D, 16'h0E5E, 16'h0E60, 16'h0E61,
16'h0E63, 16'h0E64, 16'h0E66, 16'h0E67, 16'h0E69, 16'h0E6A, 16'h0E6B, 16'h0E6D,
16'h0E6E, 16'h0E70, 16'h0E71, 16'h0E72, 16'h0E74, 16'h0E75, 16'h0E77, 16'h0E78,
16'h0E79, 16'h0E7B, 16'h0E7C, 16'h0E7E, 16'h0E7F, 16'h0E80, 16'h0E82, 16'h0E83,
16'h0E84, 16'h0E86, 16'h0E87, 16'h0E88, 16'h0E8A, 16'h0E8B, 16'h0E8C, 16'h0E8E,
16'h0E8F, 16'h0E90, 16'h0E92, 16'h0E93, 16'h0E94, 16'h0E95, 16'h0E97, 16'h0E98,
16'h0E99, 16'h0E9B, 16'h0E9C, 16'h0E9D, 16'h0E9E, 16'h0EA0, 16'h0EA1, 16'h0EA2,
16'h0EA3, 16'h0EA5, 16'h0EA6, 16'h0EA7, 16'h0EA8, 16'h0EAA, 16'h0EAB, 16'h0EAC,
16'h0EAD, 16'h0EAE, 16'h0EB0, 16'h0EB1, 16'h0EB2, 16'h0EB3, 16'h0EB4, 16'h0EB6,
16'h0EB7, 16'h0EB8, 16'h0EB9, 16'h0EBA, 16'h0EBC, 16'h0EBD, 16'h0EBE, 16'h0EBF,
16'h0EC0, 16'h0EC1, 16'h0EC2, 16'h0EC4, 16'h0EC5, 16'h0EC6, 16'h0EC7, 16'h0EC8,
16'h0EC9, 16'h0ECA, 16'h0ECC, 16'h0ECD, 16'h0ECE, 16'h0ECF, 16'h0ED0, 16'h0ED1,
16'h0ED2, 16'h0ED3, 16'h0ED4, 16'h0ED5, 16'h0ED6, 16'h0ED8, 16'h0ED9, 16'h0EDA,
16'h0EDB, 16'h0EDC, 16'h0EDD, 16'h0EDE, 16'h0EDF, 16'h0EE0, 16'h0EE1, 16'h0EE2,
16'h0EE3, 16'h0EE4, 16'h0EE5, 16'h0EE6, 16'h0EE7, 16'h0EE8, 16'h0EE9, 16'h0EEA,
16'h0EEB, 16'h0EEC, 16'h0EED, 16'h0EEE, 16'h0EEF, 16'h0EF0, 16'h0EF1, 16'h0EF2,
16'h0EF3, 16'h0EF4, 16'h0EF5, 16'h0EF6, 16'h0EF7, 16'h0EF8, 16'h0EF9, 16'h0EFA,
16'h0EFB, 16'h0EFC, 16'h0EFD, 16'h0EFE, 16'h0EFF, 16'h0F00, 16'h0F01, 16'h0F02,
16'h0F03, 16'h0F03, 16'h0F04, 16'h0F05, 16'h0F06, 16'h0F07, 16'h0F08, 16'h0F09,
16'h0F0A, 16'h0F0B, 16'h0F0C, 16'h0F0D, 16'h0F0D, 16'h0F0E, 16'h0F0F, 16'h0F10,
16'h0F11, 16'h0F12, 16'h0F13, 16'h0F14, 16'h0F15, 16'h0F15, 16'h0F16, 16'h0F17,
16'h0F18, 16'h0F19, 16'h0F1A, 16'h0F1B, 16'h0F1B, 16'h0F1C, 16'h0F1D, 16'h0F1E,
16'h0F1F, 16'h0F20, 16'h0F20, 16'h0F21, 16'h0F22, 16'h0F23, 16'h0F24, 16'h0F24,
16'h0F25, 16'h0F26, 16'h0F27, 16'h0F28, 16'h0F28, 16'h0F29, 16'h0F2A, 16'h0F2B,
16'h0F2C, 16'h0F2C, 16'h0F2D, 16'h0F2E, 16'h0F2F, 16'h0F30, 16'h0F30, 16'h0F31,
16'h0F32, 16'h0F33, 16'h0F33, 16'h0F34, 16'h0F35, 16'h0F36, 16'h0F36, 16'h0F37,
16'h0F38, 16'h0F39, 16'h0F39, 16'h0F3A, 16'h0F3B, 16'h0F3C, 16'h0F3C, 16'h0F3D,
16'h0F3E, 16'h0F3E, 16'h0F3F, 16'h0F40, 16'h0F41, 16'h0F41, 16'h0F42, 16'h0F43,
16'h0F43, 16'h0F44, 16'h0F45, 16'h0F46, 16'h0F46, 16'h0F47, 16'h0F48, 16'h0F48,
16'h0F49, 16'h0F4A, 16'h0F4A, 16'h0F4B, 16'h0F4C, 16'h0F4C, 16'h0F4D, 16'h0F4E,
16'h0F4E, 16'h0F4F, 16'h0F50, 16'h0F50, 16'h0F51, 16'h0F52, 16'h0F52, 16'h0F53,
16'h0F54, 16'h0F54, 16'h0F55, 16'h0F56, 16'h0F56, 16'h0F57, 16'h0F57, 16'h0F58,
16'h0F59, 16'h0F59, 16'h0F5A, 16'h0F5B, 16'h0F5B, 16'h0F5C, 16'h0F5C, 16'h0F5D,
16'h0F5E, 16'h0F5E, 16'h0F5F, 16'h0F5F, 16'h0F60, 16'h0F61, 16'h0F61, 16'h0F62,
16'h0F62, 16'h0F63, 16'h0F64, 16'h0F64, 16'h0F65, 16'h0F65, 16'h0F66, 16'h0F67,
16'h0F67, 16'h0F68, 16'h0F68, 16'h0F69, 16'h0F69, 16'h0F6A, 16'h0F6B, 16'h0F6B,
16'h0F6C, 16'h0F6C, 16'h0F6D, 16'h0F6D, 16'h0F6E, 16'h0F6E, 16'h0F6F, 16'h0F70,
16'h0F70, 16'h0F71, 16'h0F71, 16'h0F72, 16'h0F72, 16'h0F73, 16'h0F73, 16'h0F74,
16'h0F74, 16'h0F75, 16'h0F75, 16'h0F76, 16'h0F76, 16'h0F77, 16'h0F77, 16'h0F78,
16'h0F78, 16'h0F79, 16'h0F79, 16'h0F7A, 16'h0F7B, 16'h0F7B, 16'h0F7C, 16'h0F7C,
16'h0F7D, 16'h0F7D, 16'h0F7E, 16'h0F7E, 16'h0F7E, 16'h0F7F, 16'h0F7F, 16'h0F80,
16'h0F80, 16'h0F81, 16'h0F81, 16'h0F82, 16'h0F82, 16'h0F83, 16'h0F83, 16'h0F84,
16'h0F84, 16'h0F85, 16'h0F85, 16'h0F86, 16'h0F86, 16'h0F87, 16'h0F87, 16'h0F87,
16'h0F88, 16'h0F88, 16'h0F89, 16'h0F89, 16'h0F8A, 16'h0F8A, 16'h0F8B, 16'h0F8B,
16'h0F8C, 16'h0F8C, 16'h0F8C, 16'h0F8D, 16'h0F8D, 16'h0F8E, 16'h0F8E, 16'h0F8F,
16'h0F8F, 16'h0F8F, 16'h0F90, 16'h0F90, 16'h0F91, 16'h0F91, 16'h0F92, 16'h0F92,
16'h0F92, 16'h0F93, 16'h0F93, 16'h0F94, 16'h0F94, 16'h0F94, 16'h0F95, 16'h0F95,
16'h0F96, 16'h0F96, 16'h0F96, 16'h0F97, 16'h0F97, 16'h0F98, 16'h0F98, 16'h0F98,
16'h0F99, 16'h0F99, 16'h0F9A, 16'h0F9A, 16'h0F9A, 16'h0F9B, 16'h0F9B, 16'h0F9C,
16'h0F9C, 16'h0F9C, 16'h0F9D, 16'h0F9D, 16'h0F9D, 16'h0F9E, 16'h0F9E, 16'h0F9F,
16'h0F9F, 16'h0F9F, 16'h0FA0, 16'h0FA0, 16'h0FA0, 16'h0FA1, 16'h0FA1, 16'h0FA2,
16'h0FA2, 16'h0FA2, 16'h0FA3, 16'h0FA3, 16'h0FA3, 16'h0FA4, 16'h0FA4, 16'h0FA4,
16'h0FA5, 16'h0FA5, 16'h0FA5, 16'h0FA6, 16'h0FA6, 16'h0FA6, 16'h0FA7, 16'h0FA7,
16'h0FA7, 16'h0FA8, 16'h0FA8, 16'h0FA8, 16'h0FA9, 16'h0FA9, 16'h0FA9, 16'h0FAA,
16'h0FAA, 16'h0FAA, 16'h0FAB, 16'h0FAB, 16'h0FAB, 16'h0FAC, 16'h0FAC, 16'h0FAC,
16'h0FAD, 16'h0FAD, 16'h0FAD, 16'h0FAE, 16'h0FAE, 16'h0FAE, 16'h0FAF, 16'h0FAF,
16'h0FAF, 16'h0FB0, 16'h0FB0, 16'h0FB0, 16'h0FB0, 16'h0FB1, 16'h0FB1, 16'h0FB1,
16'h0FB2, 16'h0FB2, 16'h0FB2, 16'h0FB3, 16'h0FB3, 16'h0FB3, 16'h0FB3, 16'h0FB4,
16'h0FB4, 16'h0FB4, 16'h0FB5, 16'h0FB5, 16'h0FB5, 16'h0FB5, 16'h0FB6, 16'h0FB6,
16'h0FB6, 16'h0FB7, 16'h0FB7, 16'h0FB7, 16'h0FB7, 16'h0FB8, 16'h0FB8, 16'h0FB8,
16'h0FB9, 16'h0FB9, 16'h0FB9, 16'h0FB9, 16'h0FBA, 16'h0FBA, 16'h0FBA, 16'h0FBA,
16'h0FBB, 16'h0FBB, 16'h0FBB, 16'h0FBC, 16'h0FBC, 16'h0FBC, 16'h0FBC, 16'h0FBD,
16'h0FBD, 16'h0FBD, 16'h0FBD, 16'h0FBE, 16'h0FBE, 16'h0FBE, 16'h0FBE, 16'h0FBF,
16'h0FBF, 16'h0FBF, 16'h0FBF, 16'h0FC0, 16'h0FC0, 16'h0FC0, 16'h0FC0, 16'h0FC1,
16'h0FC1, 16'h0FC1, 16'h0FC1, 16'h0FC2, 16'h0FC2, 16'h0FC2, 16'h0FC2, 16'h0FC2,
16'h0FC3, 16'h0FC3, 16'h0FC3, 16'h0FC3, 16'h0FC4, 16'h0FC4, 16'h0FC4, 16'h0FC4,
16'h0FC5, 16'h0FC5, 16'h0FC5, 16'h0FC5, 16'h0FC6, 16'h0FC6, 16'h0FC6, 16'h0FC6,
16'h0FC6, 16'h0FC7, 16'h0FC7, 16'h0FC7, 16'h0FC7, 16'h0FC7, 16'h0FC8, 16'h0FC8,
16'h0FC8, 16'h0FC8, 16'h0FC9, 16'h0FC9, 16'h0FC9, 16'h0FC9, 16'h0FC9, 16'h0FCA,
16'h0FCA, 16'h0FCA, 16'h0FCA, 16'h0FCA, 16'h0FCB, 16'h0FCB, 16'h0FCB, 16'h0FCB,
16'h0FCB, 16'h0FCC, 16'h0FCC, 16'h0FCC, 16'h0FCC, 16'h0FCC, 16'h0FCD, 16'h0FCD,
16'h0FCD, 16'h0FCD, 16'h0FCD, 16'h0FCE, 16'h0FCE, 16'h0FCE, 16'h0FCE, 16'h0FCE,
16'h0FCF, 16'h0FCF, 16'h0FCF, 16'h0FCF, 16'h0FCF, 16'h0FD0, 16'h0FD0, 16'h0FD0,
16'h0FD0, 16'h0FD0, 16'h0FD0, 16'h0FD1, 16'h0FD1, 16'h0FD1, 16'h0FD1, 16'h0FD1,
16'h0FD2, 16'h0FD2, 16'h0FD2, 16'h0FD2, 16'h0FD2, 16'h0FD2, 16'h0FD3, 16'h0FD3,
16'h0FD3, 16'h0FD3, 16'h0FD3, 16'h0FD4, 16'h0FD4, 16'h0FD4, 16'h0FD4, 16'h0FD4,
16'h0FD4, 16'h0FD5, 16'h0FD5, 16'h0FD5, 16'h0FD5, 16'h0FD5, 16'h0FD5, 16'h0FD6,
16'h0FD6, 16'h0FD6, 16'h0FD6, 16'h0FD6, 16'h0FD6, 16'h0FD7, 16'h0FD7, 16'h0FD7,
16'h0FD7, 16'h0FD7, 16'h0FD7, 16'h0FD7, 16'h0FD8, 16'h0FD8, 16'h0FD8, 16'h0FD8,
16'h0FD8, 16'h0FD8, 16'h0FD9, 16'h0FD9, 16'h0FD9, 16'h0FD9, 16'h0FD9, 16'h0FD9,
16'h0FD9, 16'h0FDA, 16'h0FDA, 16'h0FDA, 16'h0FDA, 16'h0FDA, 16'h0FDA, 16'h0FDA,
16'h0FDB, 16'h0FDB, 16'h0FDB, 16'h0FDB, 16'h0FDB, 16'h0FDB, 16'h0FDB, 16'h0FDC,
16'h0FDC, 16'h0FDC, 16'h0FDC, 16'h0FDC, 16'h0FDC, 16'h0FDC, 16'h0FDD, 16'h0FDD,
16'h0FDD, 16'h0FDD, 16'h0FDD, 16'h0FDD, 16'h0FDD, 16'h0FDE, 16'h0FDE, 16'h0FDE,
16'h0FDE, 16'h0FDE, 16'h0FDE, 16'h0FDE, 16'h0FDE, 16'h0FDF, 16'h0FDF, 16'h0FDF,
16'h0FDF, 16'h0FDF, 16'h0FDF, 16'h0FDF, 16'h0FDF, 16'h0FE0, 16'h0FE0, 16'h0FE0,
16'h0FE0, 16'h0FE0, 16'h0FE0, 16'h0FE0, 16'h0FE0, 16'h0FE1, 16'h0FE1, 16'h0FE1,
16'h0FE1, 16'h0FE1, 16'h0FE1, 16'h0FE1, 16'h0FE1, 16'h0FE2, 16'h0FE2, 16'h0FE2,
16'h0FE2, 16'h0FE2, 16'h0FE2, 16'h0FE2, 16'h0FE2, 16'h0FE2, 16'h0FE3, 16'h0FE3,
16'h0FE3, 16'h0FE3, 16'h0FE3, 16'h0FE3, 16'h0FE3, 16'h0FE3, 16'h0FE4, 16'h0FE4,
16'h0FE4, 16'h0FE4, 16'h0FE4, 16'h0FE4, 16'h0FE4, 16'h0FE4, 16'h0FE4, 16'h0FE4,
16'h0FE5, 16'h0FE5, 16'h0FE5, 16'h0FE5, 16'h0FE5, 16'h0FE5, 16'h0FE5, 16'h0FE5,
16'h0FE5, 16'h0FE6, 16'h0FE6, 16'h0FE6, 16'h0FE6, 16'h0FE6, 16'h0FE6, 16'h0FE6,
16'h0FE6, 16'h0FE6, 16'h0FE6, 16'h0FE7, 16'h0FE7, 16'h0FE7, 16'h0FE7, 16'h0FE7,
16'h0FE7, 16'h0FE7, 16'h0FE7, 16'h0FE7, 16'h0FE7, 16'h0FE8, 16'h0FE8, 16'h0FE8,
16'h0FE8, 16'h0FE8, 16'h0FE8, 16'h0FE8, 16'h0FE8, 16'h0FE8, 16'h0FE8, 16'h0FE8,
16'h0FE9, 16'h0FE9, 16'h0FE9, 16'h0FE9, 16'h0FE9, 16'h0FE9, 16'h0FE9, 16'h0FE9,
16'h0FE9, 16'h0FE9, 16'h0FE9, 16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEA,
16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEA, 16'h0FEB,
16'h0FEB, 16'h0FEB, 16'h0FEB, 16'h0FEB, 16'h0FEB, 16'h0FEB, 16'h0FEB, 16'h0FEB,
16'h0FEB, 16'h0FEB, 16'h0FEB, 16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC,
16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC, 16'h0FEC,
16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED,
16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FED, 16'h0FEE, 16'h0FEE,
16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEE,
16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEE, 16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FEF,
16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FEF,
16'h0FEF, 16'h0FEF, 16'h0FEF, 16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0,
16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF0,
16'h0FF0, 16'h0FF0, 16'h0FF0, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1,
16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1,
16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF1, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2,
16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2,
16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF2, 16'h0FF3,
16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3,
16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3, 16'h0FF3,
16'h0FF3, 16'h0FF3, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4,
16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4,
16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4, 16'h0FF4,
16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5,
16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5,
16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF5, 16'h0FF6,
16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6,
16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6,
16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6, 16'h0FF6,
16'h0FF6, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7,
16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7,
16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7,
16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF7, 16'h0FF8, 16'h0FF8, 16'h0FF8,
16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8,
16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8,
16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8,
16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF8, 16'h0FF9, 16'h0FF9,
16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9,
16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9,
16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9,
16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9, 16'h0FF9,
16'h0FF9, 16'h0FF9, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA,
16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA,
16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA,
16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA,
16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA,
16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFA, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB, 16'h0FFB,
16'h0FFB, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC, 16'h0FFC,
16'h0FFC, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD,
16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFD, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE, 16'h0FFE,
16'h0FFE, 16'h0FFE, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h0FFF,
16'h0FFF, 16'h0FFF, 16'h0FFF, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000, 16'h1000,
16'h0800, 16'h07FC, 16'h07F8, 16'h07F4, 16'h07F0, 16'h07EC, 16'h07E8, 16'h07E4,
16'h07E0, 16'h07DC, 16'h07D8, 16'h07D4, 16'h07D0, 16'h07CC, 16'h07C8, 16'h07C4,
16'h07C0, 16'h07BC, 16'h07B8, 16'h07B4, 16'h07B0, 16'h07AC, 16'h07A8, 16'h07A4,
16'h07A0, 16'h079C, 16'h0798, 16'h0794, 16'h0790, 16'h078C, 16'h0788, 16'h0784,
16'h0780, 16'h077C, 16'h0778, 16'h0774, 16'h0770, 16'h076C, 16'h0768, 16'h0764,
16'h0760, 16'h075C, 16'h0758, 16'h0754, 16'h0750, 16'h074C, 16'h0748, 16'h0745,
16'h0741, 16'h073D, 16'h0739, 16'h0735, 16'h0731, 16'h072D, 16'h0729, 16'h0725,
16'h0721, 16'h071D, 16'h0719, 16'h0715, 16'h0711, 16'h070D, 16'h0709, 16'h0705,
16'h0701, 16'h06FD, 16'h06F9, 16'h06F6, 16'h06F2, 16'h06EE, 16'h06EA, 16'h06E6,
16'h06E2, 16'h06DE, 16'h06DA, 16'h06D6, 16'h06D2, 16'h06CE, 16'h06CA, 16'h06C6,
16'h06C3, 16'h06BF, 16'h06BB, 16'h06B7, 16'h06B3, 16'h06AF, 16'h06AB, 16'h06A7,
16'h06A3, 16'h06A0, 16'h069C, 16'h0698, 16'h0694, 16'h0690, 16'h068C, 16'h0688,
16'h0684, 16'h0681, 16'h067D, 16'h0679, 16'h0675, 16'h0671, 16'h066D, 16'h0669,
16'h0666, 16'h0662, 16'h065E, 16'h065A, 16'h0656, 16'h0652, 16'h064F, 16'h064B,
16'h0647, 16'h0643, 16'h063F, 16'h063C, 16'h0638, 16'h0634, 16'h0630, 16'h062C,
16'h0629, 16'h0625, 16'h0621, 16'h061D, 16'h0619, 16'h0616, 16'h0612, 16'h060E,
16'h060A, 16'h0607, 16'h0603, 16'h05FF, 16'h05FB, 16'h05F8, 16'h05F4, 16'h05F0,
16'h05EC, 16'h05E9, 16'h05E5, 16'h05E1, 16'h05DE, 16'h05DA, 16'h05D6, 16'h05D2,
16'h05CF, 16'h05CB, 16'h05C7, 16'h05C4, 16'h05C0, 16'h05BC, 16'h05B9, 16'h05B5,
16'h05B1, 16'h05AE, 16'h05AA, 16'h05A6, 16'h05A3, 16'h059F, 16'h059B, 16'h0598,
16'h0594, 16'h0590, 16'h058D, 16'h0589, 16'h0586, 16'h0582, 16'h057E, 16'h057B,
16'h0577, 16'h0574, 16'h0570, 16'h056C, 16'h0569, 16'h0565, 16'h0562, 16'h055E,
16'h055A, 16'h0557, 16'h0553, 16'h0550, 16'h054C, 16'h0549, 16'h0545, 16'h0542,
16'h053E, 16'h053B, 16'h0537, 16'h0534, 16'h0530, 16'h052D, 16'h0529, 16'h0526,
16'h0522, 16'h051F, 16'h051B, 16'h0518, 16'h0514, 16'h0511, 16'h050D, 16'h050A,
16'h0506, 16'h0503, 16'h04FF, 16'h04FC, 16'h04F9, 16'h04F5, 16'h04F2, 16'h04EE,
16'h04EB, 16'h04E8, 16'h04E4, 16'h04E1, 16'h04DD, 16'h04DA, 16'h04D7, 16'h04D3,
16'h04D0, 16'h04CC, 16'h04C9, 16'h04C6, 16'h04C2, 16'h04BF, 16'h04BC, 16'h04B8,
16'h04B5, 16'h04B2, 16'h04AE, 16'h04AB, 16'h04A8, 16'h04A5, 16'h04A1, 16'h049E,
16'h049B, 16'h0497, 16'h0494, 16'h0491, 16'h048E, 16'h048A, 16'h0487, 16'h0484,
16'h0481, 16'h047D, 16'h047A, 16'h0477, 16'h0474, 16'h0471, 16'h046D, 16'h046A,
16'h0467, 16'h0464, 16'h0461, 16'h045D, 16'h045A, 16'h0457, 16'h0454, 16'h0451,
16'h044E, 16'h044A, 16'h0447, 16'h0444, 16'h0441, 16'h043E, 16'h043B, 16'h0438,
16'h0435, 16'h0432, 16'h042E, 16'h042B, 16'h0428, 16'h0425, 16'h0422, 16'h041F,
16'h041C, 16'h0419, 16'h0416, 16'h0413, 16'h0410, 16'h040D, 16'h040A, 16'h0407,
16'h0404, 16'h0401, 16'h03FE, 16'h03FB, 16'h03F8, 16'h03F5, 16'h03F2, 16'h03EF,
16'h03EC, 16'h03E9, 16'h03E6, 16'h03E3, 16'h03E0, 16'h03DD, 16'h03DA, 16'h03D7,
16'h03D4, 16'h03D1, 16'h03CF, 16'h03CC, 16'h03C9, 16'h03C6, 16'h03C3, 16'h03C0,
16'h03BD, 16'h03BA, 16'h03B8, 16'h03B5, 16'h03B2, 16'h03AF, 16'h03AC, 16'h03A9,
16'h03A7, 16'h03A4, 16'h03A1, 16'h039E, 16'h039B, 16'h0399, 16'h0396, 16'h0393,
16'h0390, 16'h038D, 16'h038B, 16'h0388, 16'h0385, 16'h0382, 16'h0380, 16'h037D,
16'h037A, 16'h0377, 16'h0375, 16'h0372, 16'h036F, 16'h036D, 16'h036A, 16'h0367,
16'h0365, 16'h0362, 16'h035F, 16'h035D, 16'h035A, 16'h0357, 16'h0355, 16'h0352,
16'h034F, 16'h034D, 16'h034A, 16'h0348, 16'h0345, 16'h0342, 16'h0340, 16'h033D,
16'h033B, 16'h0338, 16'h0335, 16'h0333, 16'h0330, 16'h032E, 16'h032B, 16'h0329,
16'h0326, 16'h0324, 16'h0321, 16'h031F, 16'h031C, 16'h031A, 16'h0317, 16'h0315,
16'h0312, 16'h0310, 16'h030D, 16'h030B, 16'h0308, 16'h0306, 16'h0303, 16'h0301,
16'h02FE, 16'h02FC, 16'h02FA, 16'h02F7, 16'h02F5, 16'h02F2, 16'h02F0, 16'h02EE,
16'h02EB, 16'h02E9, 16'h02E6, 16'h02E4, 16'h02E2, 16'h02DF, 16'h02DD, 16'h02DB,
16'h02D8, 16'h02D6, 16'h02D4, 16'h02D1, 16'h02CF, 16'h02CD, 16'h02CA, 16'h02C8,
16'h02C6, 16'h02C3, 16'h02C1, 16'h02BF, 16'h02BD, 16'h02BA, 16'h02B8, 16'h02B6,
16'h02B4, 16'h02B1, 16'h02AF, 16'h02AD, 16'h02AB, 16'h02A8, 16'h02A6, 16'h02A4,
16'h02A2, 16'h02A0, 16'h029D, 16'h029B, 16'h0299, 16'h0297, 16'h0295, 16'h0293,
16'h0290, 16'h028E, 16'h028C, 16'h028A, 16'h0288, 16'h0286, 16'h0284, 16'h0282,
16'h027F, 16'h027D, 16'h027B, 16'h0279, 16'h0277, 16'h0275, 16'h0273, 16'h0271,
16'h026F, 16'h026D, 16'h026B, 16'h0269, 16'h0267, 16'h0264, 16'h0262, 16'h0260,
16'h025E, 16'h025C, 16'h025A, 16'h0258, 16'h0256, 16'h0254, 16'h0252, 16'h0250,
16'h024E, 16'h024C, 16'h024A, 16'h0249, 16'h0247, 16'h0245, 16'h0243, 16'h0241,
16'h023F, 16'h023D, 16'h023B, 16'h0239, 16'h0237, 16'h0235, 16'h0233, 16'h0231,
16'h0230, 16'h022E, 16'h022C, 16'h022A, 16'h0228, 16'h0226, 16'h0224, 16'h0222,
16'h0221, 16'h021F, 16'h021D, 16'h021B, 16'h0219, 16'h0217, 16'h0216, 16'h0214,
16'h0212, 16'h0210, 16'h020E, 16'h020D, 16'h020B, 16'h0209, 16'h0207, 16'h0206,
16'h0204, 16'h0202, 16'h0200, 16'h01FF, 16'h01FD, 16'h01FB, 16'h01F9, 16'h01F8,
16'h01F6, 16'h01F4, 16'h01F2, 16'h01F1, 16'h01EF, 16'h01ED, 16'h01EC, 16'h01EA,
16'h01E8, 16'h01E7, 16'h01E5, 16'h01E3, 16'h01E2, 16'h01E0, 16'h01DE, 16'h01DD,
16'h01DB, 16'h01D9, 16'h01D8, 16'h01D6, 16'h01D4, 16'h01D3, 16'h01D1, 16'h01D0,
16'h01CE, 16'h01CC, 16'h01CB, 16'h01C9, 16'h01C8, 16'h01C6, 16'h01C4, 16'h01C3,
16'h01C1, 16'h01C0, 16'h01BE, 16'h01BD, 16'h01BB, 16'h01BA, 16'h01B8, 16'h01B7,
16'h01B5, 16'h01B3, 16'h01B2, 16'h01B0, 16'h01AF, 16'h01AD, 16'h01AC, 16'h01AA,
16'h01A9, 16'h01A7, 16'h01A6, 16'h01A5, 16'h01A3, 16'h01A2, 16'h01A0, 16'h019F,
16'h019D, 16'h019C, 16'h019A, 16'h0199, 16'h0197, 16'h0196, 16'h0195, 16'h0193,
16'h0192, 16'h0190, 16'h018F, 16'h018E, 16'h018C, 16'h018B, 16'h0189, 16'h0188,
16'h0187, 16'h0185, 16'h0184, 16'h0182, 16'h0181, 16'h0180, 16'h017E, 16'h017D,
16'h017C, 16'h017A, 16'h0179, 16'h0178, 16'h0176, 16'h0175, 16'h0174, 16'h0172,
16'h0171, 16'h0170, 16'h016E, 16'h016D, 16'h016C, 16'h016B, 16'h0169, 16'h0168,
16'h0167, 16'h0165, 16'h0164, 16'h0163, 16'h0162, 16'h0160, 16'h015F, 16'h015E,
16'h015D, 16'h015B, 16'h015A, 16'h0159, 16'h0158, 16'h0156, 16'h0155, 16'h0154,
16'h0153, 16'h0152, 16'h0150, 16'h014F, 16'h014E, 16'h014D, 16'h014C, 16'h014A,
16'h0149, 16'h0148, 16'h0147, 16'h0146, 16'h0144, 16'h0143, 16'h0142, 16'h0141,
16'h0140, 16'h013F, 16'h013E, 16'h013C, 16'h013B, 16'h013A, 16'h0139, 16'h0138,
16'h0137, 16'h0136, 16'h0134, 16'h0133, 16'h0132, 16'h0131, 16'h0130, 16'h012F,
16'h012E, 16'h012D, 16'h012C, 16'h012B, 16'h012A, 16'h0128, 16'h0127, 16'h0126,
16'h0125, 16'h0124, 16'h0123, 16'h0122, 16'h0121, 16'h0120, 16'h011F, 16'h011E,
16'h011D, 16'h011C, 16'h011B, 16'h011A, 16'h0119, 16'h0118, 16'h0117, 16'h0116,
16'h0115, 16'h0114, 16'h0113, 16'h0112, 16'h0111, 16'h0110, 16'h010F, 16'h010E,
16'h010D, 16'h010C, 16'h010B, 16'h010A, 16'h0109, 16'h0108, 16'h0107, 16'h0106,
16'h0105, 16'h0104, 16'h0103, 16'h0102, 16'h0101, 16'h0100, 16'h00FF, 16'h00FE,
16'h00FD, 16'h00FD, 16'h00FC, 16'h00FB, 16'h00FA, 16'h00F9, 16'h00F8, 16'h00F7,
16'h00F6, 16'h00F5, 16'h00F4, 16'h00F3, 16'h00F3, 16'h00F2, 16'h00F1, 16'h00F0,
16'h00EF, 16'h00EE, 16'h00ED, 16'h00EC, 16'h00EB, 16'h00EB, 16'h00EA, 16'h00E9,
16'h00E8, 16'h00E7, 16'h00E6, 16'h00E5, 16'h00E5, 16'h00E4, 16'h00E3, 16'h00E2,
16'h00E1, 16'h00E0, 16'h00E0, 16'h00DF, 16'h00DE, 16'h00DD, 16'h00DC, 16'h00DC,
16'h00DB, 16'h00DA, 16'h00D9, 16'h00D8, 16'h00D8, 16'h00D7, 16'h00D6, 16'h00D5,
16'h00D4, 16'h00D4, 16'h00D3, 16'h00D2, 16'h00D1, 16'h00D0, 16'h00D0, 16'h00CF,
16'h00CE, 16'h00CD, 16'h00CD, 16'h00CC, 16'h00CB, 16'h00CA, 16'h00CA, 16'h00C9,
16'h00C8, 16'h00C7, 16'h00C7, 16'h00C6, 16'h00C5, 16'h00C4, 16'h00C4, 16'h00C3,
16'h00C2, 16'h00C2, 16'h00C1, 16'h00C0, 16'h00BF, 16'h00BF, 16'h00BE, 16'h00BD,
16'h00BD, 16'h00BC, 16'h00BB, 16'h00BA, 16'h00BA, 16'h00B9, 16'h00B8, 16'h00B8,
16'h00B7, 16'h00B6, 16'h00B6, 16'h00B5, 16'h00B4, 16'h00B4, 16'h00B3, 16'h00B2,
16'h00B2, 16'h00B1, 16'h00B0, 16'h00B0, 16'h00AF, 16'h00AE, 16'h00AE, 16'h00AD,
16'h00AC, 16'h00AC, 16'h00AB, 16'h00AA, 16'h00AA, 16'h00A9, 16'h00A9, 16'h00A8,
16'h00A7, 16'h00A7, 16'h00A6, 16'h00A5, 16'h00A5, 16'h00A4, 16'h00A4, 16'h00A3,
16'h00A2, 16'h00A2, 16'h00A1, 16'h00A1, 16'h00A0, 16'h009F, 16'h009F, 16'h009E,
16'h009E, 16'h009D, 16'h009C, 16'h009C, 16'h009B, 16'h009B, 16'h009A, 16'h0099,
16'h0099, 16'h0098, 16'h0098, 16'h0097, 16'h0097, 16'h0096, 16'h0095, 16'h0095,
16'h0094, 16'h0094, 16'h0093, 16'h0093, 16'h0092, 16'h0092, 16'h0091, 16'h0090,
16'h0090, 16'h008F, 16'h008F, 16'h008E, 16'h008E, 16'h008D, 16'h008D, 16'h008C,
16'h008C, 16'h008B, 16'h008B, 16'h008A, 16'h008A, 16'h0089, 16'h0089, 16'h0088,
16'h0088, 16'h0087, 16'h0087, 16'h0086, 16'h0085, 16'h0085, 16'h0084, 16'h0084,
16'h0083, 16'h0083, 16'h0082, 16'h0082, 16'h0082, 16'h0081, 16'h0081, 16'h0080,
16'h0080, 16'h007F, 16'h007F, 16'h007E, 16'h007E, 16'h007D, 16'h007D, 16'h007C,
16'h007C, 16'h007B, 16'h007B, 16'h007A, 16'h007A, 16'h0079, 16'h0079, 16'h0079,
16'h0078, 16'h0078, 16'h0077, 16'h0077, 16'h0076, 16'h0076, 16'h0075, 16'h0075,
16'h0074, 16'h0074, 16'h0074, 16'h0073, 16'h0073, 16'h0072, 16'h0072, 16'h0071,
16'h0071, 16'h0071, 16'h0070, 16'h0070, 16'h006F, 16'h006F, 16'h006E, 16'h006E,
16'h006E, 16'h006D, 16'h006D, 16'h006C, 16'h006C, 16'h006C, 16'h006B, 16'h006B,
16'h006A, 16'h006A, 16'h006A, 16'h0069, 16'h0069, 16'h0068, 16'h0068, 16'h0068,
16'h0067, 16'h0067, 16'h0066, 16'h0066, 16'h0066, 16'h0065, 16'h0065, 16'h0064,
16'h0064, 16'h0064, 16'h0063, 16'h0063, 16'h0063, 16'h0062, 16'h0062, 16'h0061,
16'h0061, 16'h0061, 16'h0060, 16'h0060, 16'h0060, 16'h005F, 16'h005F, 16'h005E,
16'h005E, 16'h005E, 16'h005D, 16'h005D, 16'h005D, 16'h005C, 16'h005C, 16'h005C,
16'h005B, 16'h005B, 16'h005B, 16'h005A, 16'h005A, 16'h005A, 16'h0059, 16'h0059,
16'h0059, 16'h0058, 16'h0058, 16'h0058, 16'h0057, 16'h0057, 16'h0057, 16'h0056,
16'h0056, 16'h0056, 16'h0055, 16'h0055, 16'h0055, 16'h0054, 16'h0054, 16'h0054,
16'h0053, 16'h0053, 16'h0053, 16'h0052, 16'h0052, 16'h0052, 16'h0051, 16'h0051,
16'h0051, 16'h0050, 16'h0050, 16'h0050, 16'h0050, 16'h004F, 16'h004F, 16'h004F,
16'h004E, 16'h004E, 16'h004E, 16'h004D, 16'h004D, 16'h004D, 16'h004D, 16'h004C,
16'h004C, 16'h004C, 16'h004B, 16'h004B, 16'h004B, 16'h004B, 16'h004A, 16'h004A,
16'h004A, 16'h0049, 16'h0049, 16'h0049, 16'h0049, 16'h0048, 16'h0048, 16'h0048,
16'h0047, 16'h0047, 16'h0047, 16'h0047, 16'h0046, 16'h0046, 16'h0046, 16'h0046,
16'h0045, 16'h0045, 16'h0045, 16'h0044, 16'h0044, 16'h0044, 16'h0044, 16'h0043,
16'h0043, 16'h0043, 16'h0043, 16'h0042, 16'h0042, 16'h0042, 16'h0042, 16'h0041,
16'h0041, 16'h0041, 16'h0041, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h003F,
16'h003F, 16'h003F, 16'h003F, 16'h003E, 16'h003E, 16'h003E, 16'h003E, 16'h003E,
16'h003D, 16'h003D, 16'h003D, 16'h003D, 16'h003C, 16'h003C, 16'h003C, 16'h003C,
16'h003B, 16'h003B, 16'h003B, 16'h003B, 16'h003A, 16'h003A, 16'h003A, 16'h003A,
16'h003A, 16'h0039, 16'h0039, 16'h0039, 16'h0039, 16'h0039, 16'h0038, 16'h0038,
16'h0038, 16'h0038, 16'h0037, 16'h0037, 16'h0037, 16'h0037, 16'h0037, 16'h0036,
16'h0036, 16'h0036, 16'h0036, 16'h0036, 16'h0035, 16'h0035, 16'h0035, 16'h0035,
16'h0035, 16'h0034, 16'h0034, 16'h0034, 16'h0034, 16'h0034, 16'h0033, 16'h0033,
16'h0033, 16'h0033, 16'h0033, 16'h0032, 16'h0032, 16'h0032, 16'h0032, 16'h0032,
16'h0031, 16'h0031, 16'h0031, 16'h0031, 16'h0031, 16'h0030, 16'h0030, 16'h0030,
16'h0030, 16'h0030, 16'h0030, 16'h002F, 16'h002F, 16'h002F, 16'h002F, 16'h002F,
16'h002E, 16'h002E, 16'h002E, 16'h002E, 16'h002E, 16'h002E, 16'h002D, 16'h002D,
16'h002D, 16'h002D, 16'h002D, 16'h002C, 16'h002C, 16'h002C, 16'h002C, 16'h002C,
16'h002C, 16'h002B, 16'h002B, 16'h002B, 16'h002B, 16'h002B, 16'h002B, 16'h002A,
16'h002A, 16'h002A, 16'h002A, 16'h002A, 16'h002A, 16'h0029, 16'h0029, 16'h0029,
16'h0029, 16'h0029, 16'h0029, 16'h0029, 16'h0028, 16'h0028, 16'h0028, 16'h0028,
16'h0028, 16'h0028, 16'h0027, 16'h0027, 16'h0027, 16'h0027, 16'h0027, 16'h0027,
16'h0027, 16'h0026, 16'h0026, 16'h0026, 16'h0026, 16'h0026, 16'h0026, 16'h0026,
16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0025, 16'h0024,
16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0024, 16'h0023, 16'h0023,
16'h0023, 16'h0023, 16'h0023, 16'h0023, 16'h0023, 16'h0022, 16'h0022, 16'h0022,
16'h0022, 16'h0022, 16'h0022, 16'h0022, 16'h0022, 16'h0021, 16'h0021, 16'h0021,
16'h0021, 16'h0021, 16'h0021, 16'h0021, 16'h0021, 16'h0020, 16'h0020, 16'h0020,
16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h0020, 16'h001F, 16'h001F, 16'h001F,
16'h001F, 16'h001F, 16'h001F, 16'h001F, 16'h001F, 16'h001E, 16'h001E, 16'h001E,
16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001E, 16'h001D, 16'h001D,
16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001D, 16'h001C, 16'h001C,
16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C, 16'h001C,
16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B, 16'h001B,
16'h001B, 16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A, 16'h001A,
16'h001A, 16'h001A, 16'h001A, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019,
16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0019, 16'h0018, 16'h0018, 16'h0018,
16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018, 16'h0018,
16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017, 16'h0017,
16'h0017, 16'h0017, 16'h0017, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016,
16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0016, 16'h0015,
16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015, 16'h0015,
16'h0015, 16'h0015, 16'h0015, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014,
16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014, 16'h0014,
16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013,
16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0013, 16'h0012, 16'h0012,
16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0012,
16'h0012, 16'h0012, 16'h0012, 16'h0012, 16'h0011, 16'h0011, 16'h0011, 16'h0011,
16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011, 16'h0011,
16'h0011, 16'h0011, 16'h0011, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010,
16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010, 16'h0010,
16'h0010, 16'h0010, 16'h0010, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F,
16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000F,
16'h000F, 16'h000F, 16'h000F, 16'h000F, 16'h000E, 16'h000E, 16'h000E, 16'h000E,
16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E,
16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000E, 16'h000D,
16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D,
16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D, 16'h000D,
16'h000D, 16'h000D, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C,
16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C,
16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C, 16'h000C,
16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B,
16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B,
16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000B, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A, 16'h000A,
16'h000A, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009,
16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0009, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008,
16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0008, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007, 16'h0007,
16'h0007, 16'h0007, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006,
16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0006, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005, 16'h0005,
16'h0005, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004, 16'h0004,
16'h0004, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003,
16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0003, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002, 16'h0002,
16'h0002, 16'h0002, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001, 16'h0001,
16'h0001, 16'h0001, 16'h0001, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000,
16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000
                                                      };
   assign out = lut[in];

endmodule // activation
