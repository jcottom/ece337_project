// $Id: $
// File name:   float_math.sv
// Created:     11/8/2016
// Author:      Cheyenne Martinez
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Floating Math Timer

module float_math
  (
    input wire start_math,
    output reg math_done
    output reg out
  );
