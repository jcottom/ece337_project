// $Id: $
// File name:   sram_buffer.sv
// Created:     11/30/2016
// Author:      Cheyenne Martinez
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: SRAM Buffer

module sram_buffer
(
	input sram_data,
	input sram_done,
	

endmodule
